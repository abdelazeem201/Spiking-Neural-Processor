/*
    ---------------------------------------------------------------------------
    Module: qspi_interface
    Author: Ahmed Abdelazeem
    Position: ASIC Design Engineer 
    ---------------------------------------------------------------------------
    Description:
        This QSPI (Quad Serial Peripheral Interface) module provides a high-speed
        interface for communication between a master device and a slave device.
        It supports full-duplex data transmission and allows for simultaneous
        reading and writing of data across multiple lines (4 data lines in this case).
        The design is intended for digital systems, such as Spiking Neural Network (SNN)
        processors, where efficient and rapid data handling is crucial.

        The QSPI interface handles data transmission in a state machine format, 
        providing functionality for both writing to and reading from the slave device
        based on the Chip Select (CS) and Serial Clock (SCK) signals.

    Parameters:
        clk        : System clock signal for synchronization.
        cs         : Chip Select signal (active low) to enable the QSPI communication.
        sck        : Serial Clock signal generated by the master device for timing.
        mosi       : Master Out Slave In data line used for sending data to the slave.
        miso       : Master In Slave Out data line used for receiving data from the slave.
        data_out   : Output register to hold the data received from the slave.

    Operation:
        - The module operates in a state machine with three states: IDLE, WRITE, and READ.
        - In the IDLE state, the module waits for the Chip Select signal to go high.
        - In the WRITE state, it captures incoming data from the MOSI line and shifts it in.
        - In the READ state, it sends the captured data out on the MISO line.
        - The transition between states is controlled by the CS signal and the SCK clock.
    ---------------------------------------------------------------------------
*/
// qspi_interface.v
module qspi_interface (
    input wire clk,               // System Clock
    input wire cs,                // Chip Select (active low)
    input wire sck,               // Serial Clock
    input wire [3:0] mosi,        // Master Out Slave In
    output reg [3:0] miso,        // Master In Slave Out
    output reg [7:0] data_out     // Data output
);
    // State definitions
    typedef enum reg [1:0] {
        IDLE = 2'b00,
        WRITE = 2'b01,
        READ = 2'b10
    } state_t;

    state_t current_state, next_state;
    reg [2:0] bit_count;           // Bit counter
    reg [7:0] data_in;            // Data input buffer

    // Sequential logic for state transition
    always @(posedge clk or negedge cs) begin
        if (!cs) begin
            current_state <= IDLE; // Reset state on Chip Select low
            bit_count <= 3'b000;    // Reset bit counter
        end else begin
            current_state <= next_state;
        end
    end

    // Combinational logic for state machine
    always @(*) begin
        next_state = current_state;
        case (current_state)
            IDLE: begin
                if (cs) begin
                    next_state = WRITE; // Move to WRITE state on CS high
                end
            end
            WRITE: begin
                if (bit_count < 3'd7) begin
                    miso <= mosi;         // Send data on MISO
                    bit_count <= bit_count + 1; // Increment bit counter
                end else begin
                    data_out <= {mosi, miso}; // Capture complete data
                    next_state = READ; // Move to READ state after write
                end
            end
            READ: begin
                if (bit_count < 3'd7) begin
                    miso <= data_out[7 - bit_count]; // Send data on MISO
                    bit_count <= bit_count + 1; // Increment bit counter
                end else begin
                    next_state = IDLE; // Return to IDLE state
                end
            end
        endcase
    end

    // Output logic for data_out and miso
    always @(posedge sck) begin
        if (current_state == WRITE) begin
            data_in <= {data_in[6:0], mosi}; // Shift in data on MOSI
        end
    end

endmodule
